`define QuickSort
//`define Matrix

`ifdef QuickSort

module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    ram_cell[       0] = 32'h000000d2;
    ram_cell[       1] = 32'h000000c3;
    ram_cell[       2] = 32'h00000099;
    ram_cell[       3] = 32'h000000a8;
    ram_cell[       4] = 32'h00000013;
    ram_cell[       5] = 32'h000000aa;
    ram_cell[       6] = 32'h00000067;
    ram_cell[       7] = 32'h00000009;
    ram_cell[       8] = 32'h00000095;
    ram_cell[       9] = 32'h00000051;
    ram_cell[      10] = 32'h000000fd;
    ram_cell[      11] = 32'h000000ab;
    ram_cell[      12] = 32'h00000014;
    ram_cell[      13] = 32'h000000d5;
    ram_cell[      14] = 32'h00000064;
    ram_cell[      15] = 32'h00000033;
    ram_cell[      16] = 32'h00000072;
    ram_cell[      17] = 32'h00000077;
    ram_cell[      18] = 32'h00000044;
    ram_cell[      19] = 32'h000000b4;
    ram_cell[      20] = 32'h0000008b;
    ram_cell[      21] = 32'h0000005d;
    ram_cell[      22] = 32'h00000001;
    ram_cell[      23] = 32'h00000045;
    ram_cell[      24] = 32'h000000f4;
    ram_cell[      25] = 32'h0000003d;
    ram_cell[      26] = 32'h00000094;
    ram_cell[      27] = 32'h000000e8;
    ram_cell[      28] = 32'h0000000f;
    ram_cell[      29] = 32'h000000d1;
    ram_cell[      30] = 32'h000000ef;
    ram_cell[      31] = 32'h00000004;
    ram_cell[      32] = 32'h000000f7;
    ram_cell[      33] = 32'h0000007f;
    ram_cell[      34] = 32'h000000f0;
    ram_cell[      35] = 32'h00000084;
    ram_cell[      36] = 32'h00000069;
    ram_cell[      37] = 32'h00000007;
    ram_cell[      38] = 32'h000000af;
    ram_cell[      39] = 32'h000000ed;
    ram_cell[      40] = 32'h00000048;
    ram_cell[      41] = 32'h000000da;
    ram_cell[      42] = 32'h00000031;
    ram_cell[      43] = 32'h00000080;
    ram_cell[      44] = 32'h000000d7;
    ram_cell[      45] = 32'h0000007d;
    ram_cell[      46] = 32'h000000c7;
    ram_cell[      47] = 32'h00000012;
    ram_cell[      48] = 32'h000000d4;
    ram_cell[      49] = 32'h0000005c;
    ram_cell[      50] = 32'h00000085;
    ram_cell[      51] = 32'h00000071;
    ram_cell[      52] = 32'h0000009d;
    ram_cell[      53] = 32'h00000027;
    ram_cell[      54] = 32'h0000006c;
    ram_cell[      55] = 32'h00000026;
    ram_cell[      56] = 32'h00000070;
    ram_cell[      57] = 32'h00000079;
    ram_cell[      58] = 32'h00000015;
    ram_cell[      59] = 32'h00000088;
    ram_cell[      60] = 32'h0000007a;
    ram_cell[      61] = 32'h000000cc;
    ram_cell[      62] = 32'h0000002e;
    ram_cell[      63] = 32'h0000004e;
    ram_cell[      64] = 32'h000000ff;
    ram_cell[      65] = 32'h0000005b;
    ram_cell[      66] = 32'h000000e4;
    ram_cell[      67] = 32'h000000f1;
    ram_cell[      68] = 32'h0000000a;
    ram_cell[      69] = 32'h0000006a;
    ram_cell[      70] = 32'h00000096;
    ram_cell[      71] = 32'h00000021;
    ram_cell[      72] = 32'h0000005e;
    ram_cell[      73] = 32'h000000bf;
    ram_cell[      74] = 32'h000000c5;
    ram_cell[      75] = 32'h000000c0;
    ram_cell[      76] = 32'h00000037;
    ram_cell[      77] = 32'h00000043;
    ram_cell[      78] = 32'h000000a2;
    ram_cell[      79] = 32'h0000000d;
    ram_cell[      80] = 32'h000000e5;
    ram_cell[      81] = 32'h00000005;
    ram_cell[      82] = 32'h00000060;
    ram_cell[      83] = 32'h0000003e;
    ram_cell[      84] = 32'h00000066;
    ram_cell[      85] = 32'h000000fb;
    ram_cell[      86] = 32'h000000dc;
    ram_cell[      87] = 32'h0000004d;
    ram_cell[      88] = 32'h00000025;
    ram_cell[      89] = 32'h000000e2;
    ram_cell[      90] = 32'h000000d0;
    ram_cell[      91] = 32'h0000002d;
    ram_cell[      92] = 32'h000000fa;
    ram_cell[      93] = 32'h00000016;
    ram_cell[      94] = 32'h0000004f;
    ram_cell[      95] = 32'h0000006f;
    ram_cell[      96] = 32'h000000ea;
    ram_cell[      97] = 32'h00000050;
    ram_cell[      98] = 32'h000000cf;
    ram_cell[      99] = 32'h00000000;
    ram_cell[     100] = 32'h000000ee;
    ram_cell[     101] = 32'h0000000b;
    ram_cell[     102] = 32'h00000040;
    ram_cell[     103] = 32'h00000059;
    ram_cell[     104] = 32'h00000054;
    ram_cell[     105] = 32'h00000082;
    ram_cell[     106] = 32'h000000de;
    ram_cell[     107] = 32'h00000055;
    ram_cell[     108] = 32'h0000002b;
    ram_cell[     109] = 32'h000000b0;
    ram_cell[     110] = 32'h00000011;
    ram_cell[     111] = 32'h0000008d;
    ram_cell[     112] = 32'h000000bb;
    ram_cell[     113] = 32'h00000098;
    ram_cell[     114] = 32'h0000009c;
    ram_cell[     115] = 32'h00000046;
    ram_cell[     116] = 32'h0000000e;
    ram_cell[     117] = 32'h000000e7;
    ram_cell[     118] = 32'h000000c4;
    ram_cell[     119] = 32'h0000009a;
    ram_cell[     120] = 32'h00000023;
    ram_cell[     121] = 32'h00000032;
    ram_cell[     122] = 32'h00000024;
    ram_cell[     123] = 32'h0000008a;
    ram_cell[     124] = 32'h000000bd;
    ram_cell[     125] = 32'h000000a0;
    ram_cell[     126] = 32'h0000008e;
    ram_cell[     127] = 32'h000000d3;
    ram_cell[     128] = 32'h00000053;
    ram_cell[     129] = 32'h0000003a;
    ram_cell[     130] = 32'h000000b1;
    ram_cell[     131] = 32'h0000009b;
    ram_cell[     132] = 32'h0000009f;
    ram_cell[     133] = 32'h000000be;
    ram_cell[     134] = 32'h000000b5;
    ram_cell[     135] = 32'h0000005a;
    ram_cell[     136] = 32'h000000e3;
    ram_cell[     137] = 32'h00000056;
    ram_cell[     138] = 32'h00000083;
    ram_cell[     139] = 32'h000000fc;
    ram_cell[     140] = 32'h000000a1;
    ram_cell[     141] = 32'h00000047;
    ram_cell[     142] = 32'h000000e6;
    ram_cell[     143] = 32'h00000074;
    ram_cell[     144] = 32'h0000001e;
    ram_cell[     145] = 32'h000000ec;
    ram_cell[     146] = 32'h000000ca;
    ram_cell[     147] = 32'h0000003b;
    ram_cell[     148] = 32'h00000028;
    ram_cell[     149] = 32'h000000fe;
    ram_cell[     150] = 32'h0000001b;
    ram_cell[     151] = 32'h00000029;
    ram_cell[     152] = 32'h00000052;
    ram_cell[     153] = 32'h00000034;
    ram_cell[     154] = 32'h00000068;
    ram_cell[     155] = 32'h00000006;
    ram_cell[     156] = 32'h0000006e;
    ram_cell[     157] = 32'h000000c9;
    ram_cell[     158] = 32'h0000008c;
    ram_cell[     159] = 32'h000000b9;
    ram_cell[     160] = 32'h000000d6;
    ram_cell[     161] = 32'h000000c8;
    ram_cell[     162] = 32'h0000002a;
    ram_cell[     163] = 32'h000000b6;
    ram_cell[     164] = 32'h0000007e;
    ram_cell[     165] = 32'h00000002;
    ram_cell[     166] = 32'h000000ae;
    ram_cell[     167] = 32'h0000003c;
    ram_cell[     168] = 32'h000000b8;
    ram_cell[     169] = 32'h00000057;
    ram_cell[     170] = 32'h0000001d;
    ram_cell[     171] = 32'h00000097;
    ram_cell[     172] = 32'h000000e0;
    ram_cell[     173] = 32'h000000bc;
    ram_cell[     174] = 32'h000000a7;
    ram_cell[     175] = 32'h00000076;
    ram_cell[     176] = 32'h00000038;
    ram_cell[     177] = 32'h000000cb;
    ram_cell[     178] = 32'h00000010;
    ram_cell[     179] = 32'h0000007c;
    ram_cell[     180] = 32'h000000ac;
    ram_cell[     181] = 32'h0000000c;
    ram_cell[     182] = 32'h000000a5;
    ram_cell[     183] = 32'h00000089;
    ram_cell[     184] = 32'h0000001f;
    ram_cell[     185] = 32'h0000006b;
    ram_cell[     186] = 32'h000000f2;
    ram_cell[     187] = 32'h0000006d;
    ram_cell[     188] = 32'h000000f8;
    ram_cell[     189] = 32'h00000036;
    ram_cell[     190] = 32'h00000042;
    ram_cell[     191] = 32'h000000c2;
    ram_cell[     192] = 32'h000000d9;
    ram_cell[     193] = 32'h00000090;
    ram_cell[     194] = 32'h00000063;
    ram_cell[     195] = 32'h000000dd;
    ram_cell[     196] = 32'h00000092;
    ram_cell[     197] = 32'h000000db;
    ram_cell[     198] = 32'h000000c6;
    ram_cell[     199] = 32'h0000009e;
    ram_cell[     200] = 32'h0000004c;
    ram_cell[     201] = 32'h000000d8;
    ram_cell[     202] = 32'h000000a6;
    ram_cell[     203] = 32'h000000ce;
    ram_cell[     204] = 32'h000000a9;
    ram_cell[     205] = 32'h000000c1;
    ram_cell[     206] = 32'h000000f3;
    ram_cell[     207] = 32'h0000001a;
    ram_cell[     208] = 32'h0000002c;
    ram_cell[     209] = 32'h00000003;
    ram_cell[     210] = 32'h00000073;
    ram_cell[     211] = 32'h00000065;
    ram_cell[     212] = 32'h0000007b;
    ram_cell[     213] = 32'h00000078;
    ram_cell[     214] = 32'h00000035;
    ram_cell[     215] = 32'h000000a3;
    ram_cell[     216] = 32'h00000087;
    ram_cell[     217] = 32'h00000022;
    ram_cell[     218] = 32'h00000061;
    ram_cell[     219] = 32'h00000017;
    ram_cell[     220] = 32'h000000f6;
    ram_cell[     221] = 32'h0000005f;
    ram_cell[     222] = 32'h0000008f;
    ram_cell[     223] = 32'h000000df;
    ram_cell[     224] = 32'h000000cd;
    ram_cell[     225] = 32'h000000b2;
    ram_cell[     226] = 32'h00000093;
    ram_cell[     227] = 32'h00000020;
    ram_cell[     228] = 32'h000000eb;
    ram_cell[     229] = 32'h00000081;
    ram_cell[     230] = 32'h00000062;
    ram_cell[     231] = 32'h000000ba;
    ram_cell[     232] = 32'h00000086;
    ram_cell[     233] = 32'h00000019;
    ram_cell[     234] = 32'h0000002f;
    ram_cell[     235] = 32'h0000001c;
    ram_cell[     236] = 32'h00000041;
    ram_cell[     237] = 32'h0000004a;
    ram_cell[     238] = 32'h000000f9;
    ram_cell[     239] = 32'h00000049;
    ram_cell[     240] = 32'h0000003f;
    ram_cell[     241] = 32'h0000004b;
    ram_cell[     242] = 32'h000000a4;
    ram_cell[     243] = 32'h000000b7;
    ram_cell[     244] = 32'h00000075;
    ram_cell[     245] = 32'h00000018;
    ram_cell[     246] = 32'h000000e1;
    ram_cell[     247] = 32'h00000058;
    ram_cell[     248] = 32'h00000039;
    ram_cell[     249] = 32'h00000030;
    ram_cell[     250] = 32'h00000008;
    ram_cell[     251] = 32'h000000f5;
    ram_cell[     252] = 32'h00000091;
    ram_cell[     253] = 32'h000000ad;
    ram_cell[     254] = 32'h000000b3;
    ram_cell[     255] = 32'h000000e9;
end

endmodule

`endif

`ifdef Matrix

module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h24212760;
    ram_cell[       1] = 32'h0;  // 32'h6af58baa;
    ram_cell[       2] = 32'h0;  // 32'h619a4d6a;
    ram_cell[       3] = 32'h0;  // 32'h6b28e2ad;
    ram_cell[       4] = 32'h0;  // 32'h365385b2;
    ram_cell[       5] = 32'h0;  // 32'ha4f8b5d5;
    ram_cell[       6] = 32'h0;  // 32'h6837ed82;
    ram_cell[       7] = 32'h0;  // 32'h2aa4dcb0;
    ram_cell[       8] = 32'h0;  // 32'hac0db735;
    ram_cell[       9] = 32'h0;  // 32'h55f7b7c3;
    ram_cell[      10] = 32'h0;  // 32'h980b2040;
    ram_cell[      11] = 32'h0;  // 32'h9b0cecf5;
    ram_cell[      12] = 32'h0;  // 32'hbf157e20;
    ram_cell[      13] = 32'h0;  // 32'h15af40e4;
    ram_cell[      14] = 32'h0;  // 32'h2edcfd50;
    ram_cell[      15] = 32'h0;  // 32'hc9c473da;
    ram_cell[      16] = 32'h0;  // 32'hdb22c107;
    ram_cell[      17] = 32'h0;  // 32'h9d388077;
    ram_cell[      18] = 32'h0;  // 32'h9328fb83;
    ram_cell[      19] = 32'h0;  // 32'h61dbb798;
    ram_cell[      20] = 32'h0;  // 32'h3d9f6055;
    ram_cell[      21] = 32'h0;  // 32'h38f33e73;
    ram_cell[      22] = 32'h0;  // 32'hd980eb25;
    ram_cell[      23] = 32'h0;  // 32'hfc2df172;
    ram_cell[      24] = 32'h0;  // 32'h844061a7;
    ram_cell[      25] = 32'h0;  // 32'hb7d7220c;
    ram_cell[      26] = 32'h0;  // 32'h3fb3694e;
    ram_cell[      27] = 32'h0;  // 32'h8b94a749;
    ram_cell[      28] = 32'h0;  // 32'h8169ce46;
    ram_cell[      29] = 32'h0;  // 32'h27d712e7;
    ram_cell[      30] = 32'h0;  // 32'h5b0cb454;
    ram_cell[      31] = 32'h0;  // 32'h3322957f;
    ram_cell[      32] = 32'h0;  // 32'h52b60a25;
    ram_cell[      33] = 32'h0;  // 32'h2658476c;
    ram_cell[      34] = 32'h0;  // 32'hd90ea95d;
    ram_cell[      35] = 32'h0;  // 32'hfd1c83f3;
    ram_cell[      36] = 32'h0;  // 32'h8ea5ba2b;
    ram_cell[      37] = 32'h0;  // 32'h0d8b9d4c;
    ram_cell[      38] = 32'h0;  // 32'h7dee1b07;
    ram_cell[      39] = 32'h0;  // 32'haf9b3288;
    ram_cell[      40] = 32'h0;  // 32'h45260b3f;
    ram_cell[      41] = 32'h0;  // 32'haa627d0b;
    ram_cell[      42] = 32'h0;  // 32'he2380f02;
    ram_cell[      43] = 32'h0;  // 32'he07da01e;
    ram_cell[      44] = 32'h0;  // 32'h3e6a6a8e;
    ram_cell[      45] = 32'h0;  // 32'he88a5546;
    ram_cell[      46] = 32'h0;  // 32'ha23d16d3;
    ram_cell[      47] = 32'h0;  // 32'hb57843be;
    ram_cell[      48] = 32'h0;  // 32'ha84ebac3;
    ram_cell[      49] = 32'h0;  // 32'hc7bc204a;
    ram_cell[      50] = 32'h0;  // 32'h6f2ba34b;
    ram_cell[      51] = 32'h0;  // 32'hb56e242d;
    ram_cell[      52] = 32'h0;  // 32'haaac9b05;
    ram_cell[      53] = 32'h0;  // 32'h29315a5a;
    ram_cell[      54] = 32'h0;  // 32'h1988ad09;
    ram_cell[      55] = 32'h0;  // 32'h98c1f0e4;
    ram_cell[      56] = 32'h0;  // 32'h8c6ea4b1;
    ram_cell[      57] = 32'h0;  // 32'h186baf86;
    ram_cell[      58] = 32'h0;  // 32'hc726866a;
    ram_cell[      59] = 32'h0;  // 32'hf8d92956;
    ram_cell[      60] = 32'h0;  // 32'h8b027e64;
    ram_cell[      61] = 32'h0;  // 32'h598055e9;
    ram_cell[      62] = 32'h0;  // 32'h2b35bf36;
    ram_cell[      63] = 32'h0;  // 32'h371d2590;
    ram_cell[      64] = 32'h0;  // 32'hcbab0c9a;
    ram_cell[      65] = 32'h0;  // 32'hff25a05f;
    ram_cell[      66] = 32'h0;  // 32'h9ff56dc6;
    ram_cell[      67] = 32'h0;  // 32'h3271b0de;
    ram_cell[      68] = 32'h0;  // 32'hf4836a16;
    ram_cell[      69] = 32'h0;  // 32'h427605cb;
    ram_cell[      70] = 32'h0;  // 32'h6a219cd2;
    ram_cell[      71] = 32'h0;  // 32'h2a8ac345;
    ram_cell[      72] = 32'h0;  // 32'h1e0865c7;
    ram_cell[      73] = 32'h0;  // 32'hb30703c1;
    ram_cell[      74] = 32'h0;  // 32'h42e89442;
    ram_cell[      75] = 32'h0;  // 32'h93e82c65;
    ram_cell[      76] = 32'h0;  // 32'hc6389e22;
    ram_cell[      77] = 32'h0;  // 32'hd080fff9;
    ram_cell[      78] = 32'h0;  // 32'h43d4ac84;
    ram_cell[      79] = 32'h0;  // 32'h178639f1;
    ram_cell[      80] = 32'h0;  // 32'h62e74ebc;
    ram_cell[      81] = 32'h0;  // 32'h66a9df43;
    ram_cell[      82] = 32'h0;  // 32'hf8f497c2;
    ram_cell[      83] = 32'h0;  // 32'hef41054a;
    ram_cell[      84] = 32'h0;  // 32'he409ced4;
    ram_cell[      85] = 32'h0;  // 32'h5d705224;
    ram_cell[      86] = 32'h0;  // 32'h09a36303;
    ram_cell[      87] = 32'h0;  // 32'h35686391;
    ram_cell[      88] = 32'h0;  // 32'h6a7bef56;
    ram_cell[      89] = 32'h0;  // 32'h0d8518b5;
    ram_cell[      90] = 32'h0;  // 32'h5b15987d;
    ram_cell[      91] = 32'h0;  // 32'ha20066dd;
    ram_cell[      92] = 32'h0;  // 32'h7710120d;
    ram_cell[      93] = 32'h0;  // 32'h25f6ffb4;
    ram_cell[      94] = 32'h0;  // 32'he8bdc551;
    ram_cell[      95] = 32'h0;  // 32'hb37cca03;
    ram_cell[      96] = 32'h0;  // 32'heefbe47c;
    ram_cell[      97] = 32'h0;  // 32'hc6bf1e9f;
    ram_cell[      98] = 32'h0;  // 32'ha675d294;
    ram_cell[      99] = 32'h0;  // 32'h36311123;
    ram_cell[     100] = 32'h0;  // 32'h8e682a73;
    ram_cell[     101] = 32'h0;  // 32'h2dba6d1b;
    ram_cell[     102] = 32'h0;  // 32'h5a631279;
    ram_cell[     103] = 32'h0;  // 32'heef3ec08;
    ram_cell[     104] = 32'h0;  // 32'h991faaae;
    ram_cell[     105] = 32'h0;  // 32'h4303c9ab;
    ram_cell[     106] = 32'h0;  // 32'h927e1329;
    ram_cell[     107] = 32'h0;  // 32'he329b743;
    ram_cell[     108] = 32'h0;  // 32'h67edbe9b;
    ram_cell[     109] = 32'h0;  // 32'hc32ff78e;
    ram_cell[     110] = 32'h0;  // 32'hd2fed818;
    ram_cell[     111] = 32'h0;  // 32'hba995387;
    ram_cell[     112] = 32'h0;  // 32'h9a05b82a;
    ram_cell[     113] = 32'h0;  // 32'hc2f94739;
    ram_cell[     114] = 32'h0;  // 32'h61855e1b;
    ram_cell[     115] = 32'h0;  // 32'h885cf825;
    ram_cell[     116] = 32'h0;  // 32'h8bdf58f0;
    ram_cell[     117] = 32'h0;  // 32'hba4e40de;
    ram_cell[     118] = 32'h0;  // 32'haacb9978;
    ram_cell[     119] = 32'h0;  // 32'he3aed9d5;
    ram_cell[     120] = 32'h0;  // 32'he3a6bdd5;
    ram_cell[     121] = 32'h0;  // 32'h9cc8ae15;
    ram_cell[     122] = 32'h0;  // 32'hc974f964;
    ram_cell[     123] = 32'h0;  // 32'h755b5822;
    ram_cell[     124] = 32'h0;  // 32'h4d9a86fc;
    ram_cell[     125] = 32'h0;  // 32'he37b06e9;
    ram_cell[     126] = 32'h0;  // 32'hdd5a0771;
    ram_cell[     127] = 32'h0;  // 32'ha698d5fb;
    ram_cell[     128] = 32'h0;  // 32'h4323a79b;
    ram_cell[     129] = 32'h0;  // 32'hffa04972;
    ram_cell[     130] = 32'h0;  // 32'h622ac7e1;
    ram_cell[     131] = 32'h0;  // 32'he0833ff0;
    ram_cell[     132] = 32'h0;  // 32'h85f543f3;
    ram_cell[     133] = 32'h0;  // 32'h52688f87;
    ram_cell[     134] = 32'h0;  // 32'h194ec7ba;
    ram_cell[     135] = 32'h0;  // 32'h6bd0adfc;
    ram_cell[     136] = 32'h0;  // 32'h053319ea;
    ram_cell[     137] = 32'h0;  // 32'h737a61f4;
    ram_cell[     138] = 32'h0;  // 32'h16176e58;
    ram_cell[     139] = 32'h0;  // 32'hf85bb8dc;
    ram_cell[     140] = 32'h0;  // 32'h85b2a446;
    ram_cell[     141] = 32'h0;  // 32'he507a79b;
    ram_cell[     142] = 32'h0;  // 32'h1d315617;
    ram_cell[     143] = 32'h0;  // 32'h36ed33c2;
    ram_cell[     144] = 32'h0;  // 32'h14bba25f;
    ram_cell[     145] = 32'h0;  // 32'hd76a55cc;
    ram_cell[     146] = 32'h0;  // 32'hc8237748;
    ram_cell[     147] = 32'h0;  // 32'hef6b32af;
    ram_cell[     148] = 32'h0;  // 32'h3e5fa6e4;
    ram_cell[     149] = 32'h0;  // 32'h52326453;
    ram_cell[     150] = 32'h0;  // 32'hac353ab0;
    ram_cell[     151] = 32'h0;  // 32'hbebb8376;
    ram_cell[     152] = 32'h0;  // 32'h5d30ba0a;
    ram_cell[     153] = 32'h0;  // 32'h9f1a1c36;
    ram_cell[     154] = 32'h0;  // 32'h7e9579b3;
    ram_cell[     155] = 32'h0;  // 32'h16844748;
    ram_cell[     156] = 32'h0;  // 32'h55beb08d;
    ram_cell[     157] = 32'h0;  // 32'h75d7f1d9;
    ram_cell[     158] = 32'h0;  // 32'hd3e3de09;
    ram_cell[     159] = 32'h0;  // 32'h466efe3e;
    ram_cell[     160] = 32'h0;  // 32'h36aa8ab1;
    ram_cell[     161] = 32'h0;  // 32'hec88e8a6;
    ram_cell[     162] = 32'h0;  // 32'h39801140;
    ram_cell[     163] = 32'h0;  // 32'had3f322b;
    ram_cell[     164] = 32'h0;  // 32'h03b3101e;
    ram_cell[     165] = 32'h0;  // 32'h71b1ecfa;
    ram_cell[     166] = 32'h0;  // 32'h1551c0a8;
    ram_cell[     167] = 32'h0;  // 32'h42c5cd12;
    ram_cell[     168] = 32'h0;  // 32'h1d3808d5;
    ram_cell[     169] = 32'h0;  // 32'haa57fe13;
    ram_cell[     170] = 32'h0;  // 32'h50194a99;
    ram_cell[     171] = 32'h0;  // 32'h48dfff90;
    ram_cell[     172] = 32'h0;  // 32'h67546bb4;
    ram_cell[     173] = 32'h0;  // 32'h9d1a2a1a;
    ram_cell[     174] = 32'h0;  // 32'h545e767c;
    ram_cell[     175] = 32'h0;  // 32'h1ae7fbb0;
    ram_cell[     176] = 32'h0;  // 32'hd416c6d6;
    ram_cell[     177] = 32'h0;  // 32'ha9f13eb8;
    ram_cell[     178] = 32'h0;  // 32'h41bb9536;
    ram_cell[     179] = 32'h0;  // 32'hd9d7a2c8;
    ram_cell[     180] = 32'h0;  // 32'hf97e2116;
    ram_cell[     181] = 32'h0;  // 32'ha65d8d46;
    ram_cell[     182] = 32'h0;  // 32'hfce94cb3;
    ram_cell[     183] = 32'h0;  // 32'h2450f5d4;
    ram_cell[     184] = 32'h0;  // 32'hac0aa5b1;
    ram_cell[     185] = 32'h0;  // 32'hc6329b2d;
    ram_cell[     186] = 32'h0;  // 32'hccd3bd94;
    ram_cell[     187] = 32'h0;  // 32'hb3b7a772;
    ram_cell[     188] = 32'h0;  // 32'h8a51ef89;
    ram_cell[     189] = 32'h0;  // 32'h704d194c;
    ram_cell[     190] = 32'h0;  // 32'h9a9d4837;
    ram_cell[     191] = 32'h0;  // 32'h95177e35;
    ram_cell[     192] = 32'h0;  // 32'h5d67956e;
    ram_cell[     193] = 32'h0;  // 32'hea21f89a;
    ram_cell[     194] = 32'h0;  // 32'hbd4d10aa;
    ram_cell[     195] = 32'h0;  // 32'h3a5d0a72;
    ram_cell[     196] = 32'h0;  // 32'hd27c0693;
    ram_cell[     197] = 32'h0;  // 32'hb2b2daba;
    ram_cell[     198] = 32'h0;  // 32'h826c8197;
    ram_cell[     199] = 32'h0;  // 32'he1f7c672;
    ram_cell[     200] = 32'h0;  // 32'h1ff69bc4;
    ram_cell[     201] = 32'h0;  // 32'hb88048d2;
    ram_cell[     202] = 32'h0;  // 32'hec896db6;
    ram_cell[     203] = 32'h0;  // 32'h47f7660a;
    ram_cell[     204] = 32'h0;  // 32'hfd8d1d97;
    ram_cell[     205] = 32'h0;  // 32'hc8aebc10;
    ram_cell[     206] = 32'h0;  // 32'habd357d7;
    ram_cell[     207] = 32'h0;  // 32'hced96ab6;
    ram_cell[     208] = 32'h0;  // 32'h97575d33;
    ram_cell[     209] = 32'h0;  // 32'hbaab9261;
    ram_cell[     210] = 32'h0;  // 32'hcb8f7eb3;
    ram_cell[     211] = 32'h0;  // 32'h3d352009;
    ram_cell[     212] = 32'h0;  // 32'h36ecda07;
    ram_cell[     213] = 32'h0;  // 32'h50d0cddd;
    ram_cell[     214] = 32'h0;  // 32'h7cda7bc6;
    ram_cell[     215] = 32'h0;  // 32'hdc87a2ea;
    ram_cell[     216] = 32'h0;  // 32'h633c182b;
    ram_cell[     217] = 32'h0;  // 32'h31a7568a;
    ram_cell[     218] = 32'h0;  // 32'hd5d967cf;
    ram_cell[     219] = 32'h0;  // 32'h27416aa6;
    ram_cell[     220] = 32'h0;  // 32'hddab5afa;
    ram_cell[     221] = 32'h0;  // 32'he53d43aa;
    ram_cell[     222] = 32'h0;  // 32'hcbd25d00;
    ram_cell[     223] = 32'h0;  // 32'h60a58b38;
    ram_cell[     224] = 32'h0;  // 32'h51680124;
    ram_cell[     225] = 32'h0;  // 32'hdf609f2c;
    ram_cell[     226] = 32'h0;  // 32'hfc4486e9;
    ram_cell[     227] = 32'h0;  // 32'h917a8a8b;
    ram_cell[     228] = 32'h0;  // 32'hdb8a96f3;
    ram_cell[     229] = 32'h0;  // 32'h35aad4e3;
    ram_cell[     230] = 32'h0;  // 32'he907ac1b;
    ram_cell[     231] = 32'h0;  // 32'h92d56fc2;
    ram_cell[     232] = 32'h0;  // 32'hc94f7b40;
    ram_cell[     233] = 32'h0;  // 32'h0782870e;
    ram_cell[     234] = 32'h0;  // 32'h22a4a27d;
    ram_cell[     235] = 32'h0;  // 32'h37cac604;
    ram_cell[     236] = 32'h0;  // 32'h29ff80ed;
    ram_cell[     237] = 32'h0;  // 32'hc77f2eca;
    ram_cell[     238] = 32'h0;  // 32'h28d6b287;
    ram_cell[     239] = 32'h0;  // 32'hc0ce4c68;
    ram_cell[     240] = 32'h0;  // 32'h34b53567;
    ram_cell[     241] = 32'h0;  // 32'h1cdf4a37;
    ram_cell[     242] = 32'h0;  // 32'h967d2bdd;
    ram_cell[     243] = 32'h0;  // 32'h39bf480f;
    ram_cell[     244] = 32'h0;  // 32'h4d3e5f6d;
    ram_cell[     245] = 32'h0;  // 32'h5048dde6;
    ram_cell[     246] = 32'h0;  // 32'h9035f183;
    ram_cell[     247] = 32'h0;  // 32'h27c16372;
    ram_cell[     248] = 32'h0;  // 32'h429b2797;
    ram_cell[     249] = 32'h0;  // 32'he05a344a;
    ram_cell[     250] = 32'h0;  // 32'h58f9b78b;
    ram_cell[     251] = 32'h0;  // 32'hda0067e3;
    ram_cell[     252] = 32'h0;  // 32'h27780ddb;
    ram_cell[     253] = 32'h0;  // 32'h7c33200d;
    ram_cell[     254] = 32'h0;  // 32'h4012dd91;
    ram_cell[     255] = 32'h0;  // 32'hf40a8020;
    // src matrix A
    ram_cell[     256] = 32'h3bbbabfc;
    ram_cell[     257] = 32'h8e6e0900;
    ram_cell[     258] = 32'h1dbe0c6d;
    ram_cell[     259] = 32'hdf443b9b;
    ram_cell[     260] = 32'hf8b86a09;
    ram_cell[     261] = 32'h9a1a340f;
    ram_cell[     262] = 32'hbbe6cdf8;
    ram_cell[     263] = 32'hdd4aabdf;
    ram_cell[     264] = 32'hde2ccc42;
    ram_cell[     265] = 32'h49b1225a;
    ram_cell[     266] = 32'h8a473646;
    ram_cell[     267] = 32'h09e206c7;
    ram_cell[     268] = 32'h845fd18b;
    ram_cell[     269] = 32'h5f76f27f;
    ram_cell[     270] = 32'h3b115850;
    ram_cell[     271] = 32'hb99a22be;
    ram_cell[     272] = 32'ha47aea33;
    ram_cell[     273] = 32'hb77bc527;
    ram_cell[     274] = 32'h17641c32;
    ram_cell[     275] = 32'h499e4f4d;
    ram_cell[     276] = 32'h35438139;
    ram_cell[     277] = 32'h142d2236;
    ram_cell[     278] = 32'h32fa3b83;
    ram_cell[     279] = 32'h38121429;
    ram_cell[     280] = 32'h90c495c6;
    ram_cell[     281] = 32'h848dad94;
    ram_cell[     282] = 32'h3e0e6966;
    ram_cell[     283] = 32'haeaf4a95;
    ram_cell[     284] = 32'h64b9e2fb;
    ram_cell[     285] = 32'hb71ffcdd;
    ram_cell[     286] = 32'hbd9bcb54;
    ram_cell[     287] = 32'h063b0c69;
    ram_cell[     288] = 32'he66fe9fe;
    ram_cell[     289] = 32'h7e7c6c51;
    ram_cell[     290] = 32'h205fb31e;
    ram_cell[     291] = 32'h2cc0e2fa;
    ram_cell[     292] = 32'hdc41a983;
    ram_cell[     293] = 32'h24e8cfa5;
    ram_cell[     294] = 32'h92a50fc9;
    ram_cell[     295] = 32'h8b77e8e8;
    ram_cell[     296] = 32'h611fa748;
    ram_cell[     297] = 32'hda911d42;
    ram_cell[     298] = 32'hf69465fd;
    ram_cell[     299] = 32'h9e565075;
    ram_cell[     300] = 32'hdd511969;
    ram_cell[     301] = 32'h1f192c25;
    ram_cell[     302] = 32'h7fbe6831;
    ram_cell[     303] = 32'hec8e5616;
    ram_cell[     304] = 32'hbdcd7000;
    ram_cell[     305] = 32'h5bcdfa17;
    ram_cell[     306] = 32'hbee32bde;
    ram_cell[     307] = 32'h3e576ba9;
    ram_cell[     308] = 32'h715a626f;
    ram_cell[     309] = 32'h2b124cea;
    ram_cell[     310] = 32'hcb34aac2;
    ram_cell[     311] = 32'he6fe5608;
    ram_cell[     312] = 32'h5a265a74;
    ram_cell[     313] = 32'h18aebce4;
    ram_cell[     314] = 32'h59dbf9be;
    ram_cell[     315] = 32'hb02e1972;
    ram_cell[     316] = 32'hb5197a4c;
    ram_cell[     317] = 32'hcec71d0e;
    ram_cell[     318] = 32'h8c87485c;
    ram_cell[     319] = 32'h2c23330d;
    ram_cell[     320] = 32'h94035479;
    ram_cell[     321] = 32'h58d12a16;
    ram_cell[     322] = 32'he7be3533;
    ram_cell[     323] = 32'hee0042c2;
    ram_cell[     324] = 32'h74b617c1;
    ram_cell[     325] = 32'h10773e89;
    ram_cell[     326] = 32'hb34e755a;
    ram_cell[     327] = 32'h591b19de;
    ram_cell[     328] = 32'h24748bc0;
    ram_cell[     329] = 32'h50569ce2;
    ram_cell[     330] = 32'h8496dd15;
    ram_cell[     331] = 32'h44bdaac6;
    ram_cell[     332] = 32'hc58bf94f;
    ram_cell[     333] = 32'h6afd1e5d;
    ram_cell[     334] = 32'h2f922e3f;
    ram_cell[     335] = 32'h9a6e80e1;
    ram_cell[     336] = 32'h15cf115c;
    ram_cell[     337] = 32'h230466a0;
    ram_cell[     338] = 32'he5ad5b37;
    ram_cell[     339] = 32'h20da2629;
    ram_cell[     340] = 32'he360f736;
    ram_cell[     341] = 32'h86d7288c;
    ram_cell[     342] = 32'h71531c33;
    ram_cell[     343] = 32'hd51c9cb9;
    ram_cell[     344] = 32'h3ec6e1cd;
    ram_cell[     345] = 32'h1c795bcb;
    ram_cell[     346] = 32'h8c607970;
    ram_cell[     347] = 32'h1cc4e0da;
    ram_cell[     348] = 32'h13c29132;
    ram_cell[     349] = 32'h395317ca;
    ram_cell[     350] = 32'h9c73ef21;
    ram_cell[     351] = 32'h95f091af;
    ram_cell[     352] = 32'h02d12b60;
    ram_cell[     353] = 32'h68dcb1df;
    ram_cell[     354] = 32'h70e37d5a;
    ram_cell[     355] = 32'h3ea39bc0;
    ram_cell[     356] = 32'he4766f13;
    ram_cell[     357] = 32'hbf0a99e5;
    ram_cell[     358] = 32'h28d4acd4;
    ram_cell[     359] = 32'h93fed28c;
    ram_cell[     360] = 32'he54e87ac;
    ram_cell[     361] = 32'h2e685c74;
    ram_cell[     362] = 32'heb79dd8e;
    ram_cell[     363] = 32'hbd1db3e3;
    ram_cell[     364] = 32'hc48ef2df;
    ram_cell[     365] = 32'hc9cc3d25;
    ram_cell[     366] = 32'hf6fcda18;
    ram_cell[     367] = 32'h006125c9;
    ram_cell[     368] = 32'h7a5a591a;
    ram_cell[     369] = 32'h333253b0;
    ram_cell[     370] = 32'h51b7de26;
    ram_cell[     371] = 32'h4a455a07;
    ram_cell[     372] = 32'hfcdedb57;
    ram_cell[     373] = 32'h045b1777;
    ram_cell[     374] = 32'h1694ffe6;
    ram_cell[     375] = 32'hfb98a586;
    ram_cell[     376] = 32'h41700d50;
    ram_cell[     377] = 32'hbef4585b;
    ram_cell[     378] = 32'hddaf74c5;
    ram_cell[     379] = 32'heb1b3fb4;
    ram_cell[     380] = 32'h06544919;
    ram_cell[     381] = 32'h4788c0dc;
    ram_cell[     382] = 32'h14f39349;
    ram_cell[     383] = 32'hb3ef94e0;
    ram_cell[     384] = 32'hae343ad4;
    ram_cell[     385] = 32'hf49b5c4e;
    ram_cell[     386] = 32'h831a8bbb;
    ram_cell[     387] = 32'hcbb7928f;
    ram_cell[     388] = 32'h4aa6d5d6;
    ram_cell[     389] = 32'h886f1d4d;
    ram_cell[     390] = 32'h4121b2f8;
    ram_cell[     391] = 32'hfee25921;
    ram_cell[     392] = 32'hf3f438dd;
    ram_cell[     393] = 32'hc41d22b1;
    ram_cell[     394] = 32'h42f3580e;
    ram_cell[     395] = 32'hf64dace1;
    ram_cell[     396] = 32'h94fcc589;
    ram_cell[     397] = 32'h2f6660ab;
    ram_cell[     398] = 32'h39d492ae;
    ram_cell[     399] = 32'hfff35645;
    ram_cell[     400] = 32'ha4083d57;
    ram_cell[     401] = 32'hd08ddb1f;
    ram_cell[     402] = 32'h0d0ed119;
    ram_cell[     403] = 32'hd10a7039;
    ram_cell[     404] = 32'h3e9cc865;
    ram_cell[     405] = 32'h9401c9b3;
    ram_cell[     406] = 32'hddbdaef3;
    ram_cell[     407] = 32'hb6bf39d1;
    ram_cell[     408] = 32'h0e0d7c89;
    ram_cell[     409] = 32'h5bbb66fa;
    ram_cell[     410] = 32'h76fcea0a;
    ram_cell[     411] = 32'hf61fead3;
    ram_cell[     412] = 32'ha3b2f7fd;
    ram_cell[     413] = 32'hfc3509db;
    ram_cell[     414] = 32'h0705e1e9;
    ram_cell[     415] = 32'hcdb45a56;
    ram_cell[     416] = 32'hfac40949;
    ram_cell[     417] = 32'hf402872e;
    ram_cell[     418] = 32'hdbecbc9a;
    ram_cell[     419] = 32'hb6172d98;
    ram_cell[     420] = 32'h31985d45;
    ram_cell[     421] = 32'ha360278d;
    ram_cell[     422] = 32'h18637bcc;
    ram_cell[     423] = 32'hcbd7be9a;
    ram_cell[     424] = 32'h33934214;
    ram_cell[     425] = 32'he1381eed;
    ram_cell[     426] = 32'h964cda50;
    ram_cell[     427] = 32'hfeb8fa2e;
    ram_cell[     428] = 32'h573bdbbe;
    ram_cell[     429] = 32'h132b66a7;
    ram_cell[     430] = 32'hb448025b;
    ram_cell[     431] = 32'h8c3c20f7;
    ram_cell[     432] = 32'ha02c70a4;
    ram_cell[     433] = 32'h19ecde50;
    ram_cell[     434] = 32'h21c6a5fd;
    ram_cell[     435] = 32'h2012f0d3;
    ram_cell[     436] = 32'h9083041e;
    ram_cell[     437] = 32'hda97adea;
    ram_cell[     438] = 32'h6e27f115;
    ram_cell[     439] = 32'h1b9766e4;
    ram_cell[     440] = 32'hb630262f;
    ram_cell[     441] = 32'h3320a94f;
    ram_cell[     442] = 32'h8fb4b2c1;
    ram_cell[     443] = 32'h7a42e0e8;
    ram_cell[     444] = 32'h1dc1a424;
    ram_cell[     445] = 32'h1db723e5;
    ram_cell[     446] = 32'h958ba05a;
    ram_cell[     447] = 32'h54d29b7c;
    ram_cell[     448] = 32'h2915e40e;
    ram_cell[     449] = 32'h9e4428de;
    ram_cell[     450] = 32'h269aedc6;
    ram_cell[     451] = 32'h1bb97193;
    ram_cell[     452] = 32'hab7dec63;
    ram_cell[     453] = 32'ha36b599d;
    ram_cell[     454] = 32'h4a5e69ac;
    ram_cell[     455] = 32'h30a25734;
    ram_cell[     456] = 32'h9b8bdd76;
    ram_cell[     457] = 32'h9cb2d401;
    ram_cell[     458] = 32'h2ef86397;
    ram_cell[     459] = 32'h0b295ff0;
    ram_cell[     460] = 32'h970de362;
    ram_cell[     461] = 32'hc4565522;
    ram_cell[     462] = 32'h1469bc46;
    ram_cell[     463] = 32'he4ec41cd;
    ram_cell[     464] = 32'hfcce8b73;
    ram_cell[     465] = 32'h40c69fb2;
    ram_cell[     466] = 32'h3619369d;
    ram_cell[     467] = 32'h183a4e24;
    ram_cell[     468] = 32'h1217fd26;
    ram_cell[     469] = 32'hea8738c8;
    ram_cell[     470] = 32'h62d33c42;
    ram_cell[     471] = 32'h87efbf00;
    ram_cell[     472] = 32'h38e75ece;
    ram_cell[     473] = 32'hefbe8b20;
    ram_cell[     474] = 32'he9df9ccb;
    ram_cell[     475] = 32'h7af3d749;
    ram_cell[     476] = 32'he3932a44;
    ram_cell[     477] = 32'h50cf6275;
    ram_cell[     478] = 32'h7a33a782;
    ram_cell[     479] = 32'hc6387f73;
    ram_cell[     480] = 32'h50d42208;
    ram_cell[     481] = 32'hd9f37a7e;
    ram_cell[     482] = 32'heb467a8e;
    ram_cell[     483] = 32'hbc20b9f5;
    ram_cell[     484] = 32'h253c05c0;
    ram_cell[     485] = 32'h644633f6;
    ram_cell[     486] = 32'hf7a47924;
    ram_cell[     487] = 32'h6856d210;
    ram_cell[     488] = 32'hb668c66f;
    ram_cell[     489] = 32'h8cad5e5f;
    ram_cell[     490] = 32'h3933ee66;
    ram_cell[     491] = 32'h61dee86b;
    ram_cell[     492] = 32'h66ca5798;
    ram_cell[     493] = 32'hce291eda;
    ram_cell[     494] = 32'hdfd7dec0;
    ram_cell[     495] = 32'h10a4edf5;
    ram_cell[     496] = 32'he0f8c78b;
    ram_cell[     497] = 32'ha26489f2;
    ram_cell[     498] = 32'h5271adaf;
    ram_cell[     499] = 32'heac3ffef;
    ram_cell[     500] = 32'h4c0d162e;
    ram_cell[     501] = 32'h7f79770c;
    ram_cell[     502] = 32'h87ec9286;
    ram_cell[     503] = 32'hf03b6d82;
    ram_cell[     504] = 32'hd43af503;
    ram_cell[     505] = 32'hd3ba6f8b;
    ram_cell[     506] = 32'ha5e37003;
    ram_cell[     507] = 32'hd2ecf919;
    ram_cell[     508] = 32'he9e6ebd0;
    ram_cell[     509] = 32'h2bfbf6ef;
    ram_cell[     510] = 32'h4ff0a54f;
    ram_cell[     511] = 32'hdb24f33f;
    // src matrix B
    ram_cell[     512] = 32'hc3746e85;
    ram_cell[     513] = 32'hfb2939e8;
    ram_cell[     514] = 32'hbc2cd0fd;
    ram_cell[     515] = 32'he6ef5f57;
    ram_cell[     516] = 32'h94d152de;
    ram_cell[     517] = 32'h77a35ec6;
    ram_cell[     518] = 32'h63f68caf;
    ram_cell[     519] = 32'h774becc0;
    ram_cell[     520] = 32'h196667db;
    ram_cell[     521] = 32'ha052662f;
    ram_cell[     522] = 32'h23345815;
    ram_cell[     523] = 32'hc0ab0dca;
    ram_cell[     524] = 32'h741fb962;
    ram_cell[     525] = 32'hf3c4dbc6;
    ram_cell[     526] = 32'h0edba6e1;
    ram_cell[     527] = 32'h6a3ec57b;
    ram_cell[     528] = 32'h0901c234;
    ram_cell[     529] = 32'hc198a8cc;
    ram_cell[     530] = 32'h19b2e2f1;
    ram_cell[     531] = 32'hc3b81f12;
    ram_cell[     532] = 32'hc757c46c;
    ram_cell[     533] = 32'h072d9f86;
    ram_cell[     534] = 32'h7d10f516;
    ram_cell[     535] = 32'h4a3669a2;
    ram_cell[     536] = 32'h28c5461c;
    ram_cell[     537] = 32'h21b8a4a2;
    ram_cell[     538] = 32'h72e0bab9;
    ram_cell[     539] = 32'h48bd186f;
    ram_cell[     540] = 32'h7619f619;
    ram_cell[     541] = 32'hadc1f6db;
    ram_cell[     542] = 32'h9201af6b;
    ram_cell[     543] = 32'h5fc6cace;
    ram_cell[     544] = 32'h31675f24;
    ram_cell[     545] = 32'hc53a9534;
    ram_cell[     546] = 32'hbce65094;
    ram_cell[     547] = 32'h2d2f07b0;
    ram_cell[     548] = 32'h9c6f7e06;
    ram_cell[     549] = 32'h47e12b3c;
    ram_cell[     550] = 32'ha71f4bc3;
    ram_cell[     551] = 32'h4c1facdd;
    ram_cell[     552] = 32'h5b29f348;
    ram_cell[     553] = 32'hb44e2288;
    ram_cell[     554] = 32'hda59b619;
    ram_cell[     555] = 32'hadbe7a28;
    ram_cell[     556] = 32'h930fd807;
    ram_cell[     557] = 32'h6a52d173;
    ram_cell[     558] = 32'hb03ef567;
    ram_cell[     559] = 32'hecaa8aee;
    ram_cell[     560] = 32'hcd0a935e;
    ram_cell[     561] = 32'hfe7088ff;
    ram_cell[     562] = 32'hb17ad512;
    ram_cell[     563] = 32'h7c632b25;
    ram_cell[     564] = 32'h69d18a45;
    ram_cell[     565] = 32'hf6a9fa73;
    ram_cell[     566] = 32'hbabdcfd8;
    ram_cell[     567] = 32'h99c8576f;
    ram_cell[     568] = 32'hf5164780;
    ram_cell[     569] = 32'he77473e1;
    ram_cell[     570] = 32'h325633e2;
    ram_cell[     571] = 32'haace9e37;
    ram_cell[     572] = 32'he1aa6f70;
    ram_cell[     573] = 32'h86de3b3e;
    ram_cell[     574] = 32'h5927e626;
    ram_cell[     575] = 32'h04b4fa2e;
    ram_cell[     576] = 32'h380f1030;
    ram_cell[     577] = 32'haff5ebf5;
    ram_cell[     578] = 32'h02f4b671;
    ram_cell[     579] = 32'h8735b8af;
    ram_cell[     580] = 32'hbc3c7a2e;
    ram_cell[     581] = 32'hdd87aaf0;
    ram_cell[     582] = 32'hfd118605;
    ram_cell[     583] = 32'hbd96072a;
    ram_cell[     584] = 32'h2670733f;
    ram_cell[     585] = 32'h195f0f67;
    ram_cell[     586] = 32'hd6986279;
    ram_cell[     587] = 32'h1331eb4b;
    ram_cell[     588] = 32'h34703549;
    ram_cell[     589] = 32'hf53a6a70;
    ram_cell[     590] = 32'h16c7050a;
    ram_cell[     591] = 32'hb75810e6;
    ram_cell[     592] = 32'he3cc44db;
    ram_cell[     593] = 32'h460d235a;
    ram_cell[     594] = 32'h719b9687;
    ram_cell[     595] = 32'h3a66969e;
    ram_cell[     596] = 32'h2e923f03;
    ram_cell[     597] = 32'h14fdfa81;
    ram_cell[     598] = 32'hd2f57f54;
    ram_cell[     599] = 32'hc2b2604c;
    ram_cell[     600] = 32'h304cdbc6;
    ram_cell[     601] = 32'ha3b91f74;
    ram_cell[     602] = 32'h73d683d0;
    ram_cell[     603] = 32'hc4273100;
    ram_cell[     604] = 32'haad83194;
    ram_cell[     605] = 32'h3cf415ab;
    ram_cell[     606] = 32'hd3c67979;
    ram_cell[     607] = 32'h65c93e1c;
    ram_cell[     608] = 32'h4e053f6a;
    ram_cell[     609] = 32'h88282cdd;
    ram_cell[     610] = 32'h4251db45;
    ram_cell[     611] = 32'h638fc7f5;
    ram_cell[     612] = 32'h30592022;
    ram_cell[     613] = 32'ha842ce9e;
    ram_cell[     614] = 32'hbd8d5f67;
    ram_cell[     615] = 32'hfa50c2ec;
    ram_cell[     616] = 32'h1456836d;
    ram_cell[     617] = 32'h96ff9a30;
    ram_cell[     618] = 32'h78e51897;
    ram_cell[     619] = 32'he335a3ae;
    ram_cell[     620] = 32'hd54a8754;
    ram_cell[     621] = 32'hb59f8834;
    ram_cell[     622] = 32'hc8ec8271;
    ram_cell[     623] = 32'h23cb854c;
    ram_cell[     624] = 32'ha0eb0bd5;
    ram_cell[     625] = 32'hb98b0da0;
    ram_cell[     626] = 32'hf6f7799a;
    ram_cell[     627] = 32'h41db3f7c;
    ram_cell[     628] = 32'h7def07be;
    ram_cell[     629] = 32'ha21a4ac2;
    ram_cell[     630] = 32'h3795f896;
    ram_cell[     631] = 32'h6ffa87eb;
    ram_cell[     632] = 32'hba5bc4eb;
    ram_cell[     633] = 32'h700a7e5b;
    ram_cell[     634] = 32'h952d2007;
    ram_cell[     635] = 32'he79883bf;
    ram_cell[     636] = 32'h2df35c33;
    ram_cell[     637] = 32'he59c2db4;
    ram_cell[     638] = 32'h9d0af229;
    ram_cell[     639] = 32'haf048cfd;
    ram_cell[     640] = 32'hcfecbae8;
    ram_cell[     641] = 32'h4b0a101d;
    ram_cell[     642] = 32'he41e92b6;
    ram_cell[     643] = 32'h03556bd4;
    ram_cell[     644] = 32'h8590f58c;
    ram_cell[     645] = 32'h5ae2b049;
    ram_cell[     646] = 32'h19b6bb1c;
    ram_cell[     647] = 32'h4f102a42;
    ram_cell[     648] = 32'h378a02bf;
    ram_cell[     649] = 32'h552373fb;
    ram_cell[     650] = 32'h3d756d95;
    ram_cell[     651] = 32'hfe3e47d3;
    ram_cell[     652] = 32'h9f81f11c;
    ram_cell[     653] = 32'hfc414c4e;
    ram_cell[     654] = 32'h437821b3;
    ram_cell[     655] = 32'h2ed62e61;
    ram_cell[     656] = 32'h0942b512;
    ram_cell[     657] = 32'h7722b002;
    ram_cell[     658] = 32'hefa1f25d;
    ram_cell[     659] = 32'h90cb7f0d;
    ram_cell[     660] = 32'h7444fca9;
    ram_cell[     661] = 32'hb7da0976;
    ram_cell[     662] = 32'hf16883a9;
    ram_cell[     663] = 32'hdc67bc61;
    ram_cell[     664] = 32'h0f568eef;
    ram_cell[     665] = 32'hbdd4a70b;
    ram_cell[     666] = 32'h68bc4e1e;
    ram_cell[     667] = 32'h0c99e348;
    ram_cell[     668] = 32'hff8337a7;
    ram_cell[     669] = 32'h5632b843;
    ram_cell[     670] = 32'hed81aae1;
    ram_cell[     671] = 32'h77fa3af9;
    ram_cell[     672] = 32'h798b9ff8;
    ram_cell[     673] = 32'ha8e2e2c2;
    ram_cell[     674] = 32'h0e81dfd8;
    ram_cell[     675] = 32'h3cab241c;
    ram_cell[     676] = 32'h378c319a;
    ram_cell[     677] = 32'h69198e4d;
    ram_cell[     678] = 32'h2ab8aced;
    ram_cell[     679] = 32'haea9714d;
    ram_cell[     680] = 32'ha299406c;
    ram_cell[     681] = 32'h91978a99;
    ram_cell[     682] = 32'h86052b3b;
    ram_cell[     683] = 32'he832994f;
    ram_cell[     684] = 32'h1fe2e363;
    ram_cell[     685] = 32'h93f24d56;
    ram_cell[     686] = 32'h47701f96;
    ram_cell[     687] = 32'h468f1e97;
    ram_cell[     688] = 32'h8530a6db;
    ram_cell[     689] = 32'hbf59b27c;
    ram_cell[     690] = 32'h5364915f;
    ram_cell[     691] = 32'hbdb38050;
    ram_cell[     692] = 32'h1a2294af;
    ram_cell[     693] = 32'h97699be4;
    ram_cell[     694] = 32'hcf37d51e;
    ram_cell[     695] = 32'h256cb6dd;
    ram_cell[     696] = 32'h1a509fae;
    ram_cell[     697] = 32'he3801ab1;
    ram_cell[     698] = 32'h00a7d050;
    ram_cell[     699] = 32'hd61fa8a5;
    ram_cell[     700] = 32'hcda04400;
    ram_cell[     701] = 32'h48292b11;
    ram_cell[     702] = 32'hfa680c96;
    ram_cell[     703] = 32'hea0dfdda;
    ram_cell[     704] = 32'h4b95d603;
    ram_cell[     705] = 32'h11677c0b;
    ram_cell[     706] = 32'hf269690d;
    ram_cell[     707] = 32'ha6a50f38;
    ram_cell[     708] = 32'hb4734621;
    ram_cell[     709] = 32'h8ada7ad6;
    ram_cell[     710] = 32'hfc7a3efd;
    ram_cell[     711] = 32'hb460be52;
    ram_cell[     712] = 32'ha0832205;
    ram_cell[     713] = 32'h00e69e40;
    ram_cell[     714] = 32'hb2312305;
    ram_cell[     715] = 32'h01629b60;
    ram_cell[     716] = 32'h57a921d1;
    ram_cell[     717] = 32'hac412fc9;
    ram_cell[     718] = 32'h5632ef16;
    ram_cell[     719] = 32'h8b2bd57d;
    ram_cell[     720] = 32'h5b7ce444;
    ram_cell[     721] = 32'h32e5ad8d;
    ram_cell[     722] = 32'h582a91e8;
    ram_cell[     723] = 32'haa92ef2d;
    ram_cell[     724] = 32'he49640a4;
    ram_cell[     725] = 32'h5dae1e09;
    ram_cell[     726] = 32'h177b4d4d;
    ram_cell[     727] = 32'h67124f56;
    ram_cell[     728] = 32'h564de21e;
    ram_cell[     729] = 32'h42bb33a1;
    ram_cell[     730] = 32'h5e50c2b0;
    ram_cell[     731] = 32'h6e2df8fb;
    ram_cell[     732] = 32'h25a076c6;
    ram_cell[     733] = 32'h74647674;
    ram_cell[     734] = 32'h9da0d553;
    ram_cell[     735] = 32'h93c20a66;
    ram_cell[     736] = 32'h1e906880;
    ram_cell[     737] = 32'hfd6fd982;
    ram_cell[     738] = 32'h42b62a03;
    ram_cell[     739] = 32'hc33082ac;
    ram_cell[     740] = 32'he6d9135c;
    ram_cell[     741] = 32'h033c457b;
    ram_cell[     742] = 32'h44a7a772;
    ram_cell[     743] = 32'h15007656;
    ram_cell[     744] = 32'h578d90ba;
    ram_cell[     745] = 32'h42ba6b17;
    ram_cell[     746] = 32'h64751ded;
    ram_cell[     747] = 32'h7b35a069;
    ram_cell[     748] = 32'h7cabe984;
    ram_cell[     749] = 32'h3d0bc2f2;
    ram_cell[     750] = 32'h206d8d49;
    ram_cell[     751] = 32'h6675495a;
    ram_cell[     752] = 32'he0c31fbb;
    ram_cell[     753] = 32'hdc14b500;
    ram_cell[     754] = 32'hd8b70425;
    ram_cell[     755] = 32'hbc931055;
    ram_cell[     756] = 32'h33d9f602;
    ram_cell[     757] = 32'h3b46d703;
    ram_cell[     758] = 32'h3e8f6d8a;
    ram_cell[     759] = 32'h4a332e9f;
    ram_cell[     760] = 32'h7711600e;
    ram_cell[     761] = 32'hbbef3080;
    ram_cell[     762] = 32'hb5da5b74;
    ram_cell[     763] = 32'h0dfe60d3;
    ram_cell[     764] = 32'h21e91c30;
    ram_cell[     765] = 32'h92ed67be;
    ram_cell[     766] = 32'hd934475d;
    ram_cell[     767] = 32'h56f9ccdc;
end

endmodule

`endif