`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: USTC ESLAB
// Engineer: Huang Yifan (hyf15@mail.ustc.edu.cn)
// 
// Design Name: RV32I Core
// Module Name: RV32I Core
// Tool Versions: Vivado 2017.4.1
// Description: Top level of our CPU Core
//////////////////////////////////////////////////////////////////////////////////


//功能说明
    // RV32I Core的顶层模块

`include "Parameters.v" 
module RV32ICore(
    input wire CPU_CLK,
    input wire CPU_RST,
    input wire [31:0] CPU_Debug_DataCache_A2,
    input wire [31:0] CPU_Debug_DataCache_WD2,
    input wire [3:0] CPU_Debug_DataCache_WE2,
    output wire [31:0] CPU_Debug_DataCache_RD2,
    input wire [31:0] CPU_Debug_InstCache_A2,
    input wire [31:0] CPU_Debug_InstCache_WD2,
    input wire [ 3:0] CPU_Debug_InstCache_WE2,
    output wire [31:0] CPU_Debug_InstCache_RD2,
    //Lab3
    output wire debug_miss,
    output wire debug_cache_hit,
    output wire [31:0]total_count,
    //Lab4
    reg [31:0] br_count,
    reg [31:0] prediction_wrong_count
    );

	//wire values definitions
    wire bubbleF, flushF, bubbleD, flushD, bubbleE, flushE, bubbleM, flushM, bubbleW, flushW;
    wire [31:0] jal_target, br_target;
    wire jal, br;
    wire jalr_ID, jalr_EX;
    wire [31:0] NPC, PC_IF, PC_4, PC_ID, PC_EX;
    wire [31:0] inst_ID;
    wire reg_write_en_ID, reg_write_en_EX, reg_write_en_MEM, reg_write_en_WB;
    wire [4:0] reg1_src_EX;
    wire [4:0] reg2_src_EX;
    wire [4:0] reg_dest_EX, reg_dest_MEM, reg_dest_WB;
    wire [31:0] data_WB;
    wire [31:0] reg1, reg1_EX;
    wire [31:0] reg2, reg2_EX, reg2_MEM;
    wire [31:0] op2;
    wire [31:0] reg_or_imm;
    wire op2_src;
    wire [3:0] ALU_func_ID, ALU_func_EX;
    wire [2:0] br_type_ID, br_type_EX;
    wire load_npc_ID, load_npc_EX;
    wire wb_select_ID, wb_select_EX, wb_select_MEM;
    wire [2:0] load_type_ID, load_type_EX, load_type_MEM;
    wire [1:0] src_reg_en_ID, src_reg_en_EX;
    wire [3:0] cache_write_en_ID, cache_write_en_EX, cache_write_en_MEM;
    wire alu_src1_ID, alu_src1_EX;
    wire [1:0] alu_src2_ID, alu_src2_EX;
    wire [2:0] imm_type;
    wire [31:0] imm;
    wire [31:0] ALU_op1, ALU_op2, ALU_out;
    wire [31:0] dealt_reg2;
    wire [31:0] result, result_MEM;
    wire [1:0] op1_sel, op2_sel, reg2_sel;

    //TODO: CSR debug
    wire [11:0] csr_addr_EX;
    wire [2:0] csr_funct3_out;
    wire [4:0] csr_zimm_out;
    wire csr_write_en_in,csr_write_en_out;
    assign csr_write_en_in = inst_ID[6:0] == `CSR ? (inst_ID[19:15] == 5'b0 ? 1'b0 :1'b1) : 1'b0;
    wire is_csr_in,is_csr_out;
    assign is_csr_in = inst_ID[6:0] == `CSR ? 1'b1 : 1'b0;
    wire [31:0] csr_read_data;


    //Lab4
    wire btb_if, btb_id, btb_ex;
    wire [31:0] prediction_if, prediction_id, prediction_ex;
    wire if_prediction_true;
    wire [1:0] btb_operation;
    
    btb_id_seg my_btb_id_seg(
        .clk(CPU_CLK),
        .bubbleD(bubbleD),
        .flushD(flushD),
        .btb_if(btb_if),
        .btb_id(btb_id),
        .prediction_if(prediction_if),
        .prediction_id(prediction_id)
    );
    
    btb_ex_seg my_btb_ex_seg(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .btb_ex(btb_ex),
        .btb_id(btb_id),
        .prediction_id(prediction_id),
        .prediction_ex(prediction_ex)
    );
    
    branch_target_buffer 
    #(
        .BUFFER_ADDR_LEN(7)
    )
    my_btb
    (
        .clk(CPU_CLK), 
        .rst(CPU_RST),
        .hit(btb_if),         
        .raddr(PC_IF+4),
        .rd_data(prediction_if),                 //Predicted target     
        .operation_type(btb_operation),          //btb operation
        .waddr(PC_EX),                           //PCE(Update addr)
        .wr_data(br_target)                      //BrcPC
    );
    
    wire bht_if, bht_id, bht_ex;
    wire [31:0] final_prediction_if, final_prediction_id, final_prediction_ex;
    assign final_prediction_if = bht_if ? (btb_if ? prediction_if : PC_IF + 8) : (PC_IF + 8);
    assign if_prediction_true = (final_prediction_ex == br_target) ? 1'b1 : 1'b0;
    assign btb_operation = br ? (btb_ex ? (if_prediction_true ? `BTB_NONE : `BTB_UPDATE) : `BTB_ADD) : (btb_ex ? ( bht_ex? `BTB_NONE:`BTB_REMOVE) : `BTB_NONE);
    
    //Lab4 test 
    initial
    begin
        br_count = 0;
        prediction_wrong_count = 0;
    end
    always@(posedge CPU_CLK or posedge CPU_RST)
    begin
    if(CPU_RST)
        begin
            br_count = 0;
            prediction_wrong_count = 0;
        end
    else
        begin
        if(inst_ID[6:0] == `BRANCH)
            begin
                br_count = br_count + 1;
            end
        if(!if_prediction_true && br || ~br && (btb_ex && bht_ex))
            begin
                prediction_wrong_count = prediction_wrong_count + 1;
            end
        end
    end
    
    localparam  bht_addr_len = 7;
    bht #(
     .BHT_ADDR_LEN(bht_addr_len)
    ) my_bht
    (
        .clk(CPU_CLK), 
        .rst(CPU_RST),
        .br_ex(br),        
        .raddr(prediction_if[bht_addr_len-1:0]),     
        .waddr(prediction_ex[bht_addr_len-1:0]),  
        .prediction_taken(bht_if)      
    );

    bht_ex_seg my_hbt_ex_seg(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .bht_id(bht_id),
        .final_prediction_id(final_prediction_id),
        .bht_ex(bht_ex),
        .final_prediction_ex(final_prediction_ex)
    );

    bht_id_seg my_hbt_id_seg(
        .clk(CPU_CLK),
        .bubbleD(bubbleD),
        .flushD(flushD),
        .bht_id(bht_id),
        .final_prediction_id(final_prediction_id),
        .bht_if(bht_if),
        .final_prediction_if(final_prediction_if)
    );
    
    // Adder to compute PC + 4
    assign PC_4 = PC_IF + 4;
    // MUX for op2 source
    assign op2 = op2_src ? imm : reg2;
    // Adder to compute PC_ID + Imm - 4
    assign jal_target = PC_ID + op2 - 4;
    // MUX for ALU op1
    assign ALU_op1 = (op1_sel == 2'h0) ? result_MEM :
                                         ((op1_sel == 2'h1) ? data_WB :
                                                              (op1_sel == 2'h2) ? (PC_EX - 4) :
                                                                                  reg1_EX);
    // MUX for ALU op2
    assign ALU_op2 = (op2_sel == 2'h0) ? result_MEM :
                                         ((op2_sel == 2'h1) ? data_WB :
                                                              ((op2_sel == 2'h2) ? reg2_src_EX :
                                                                                   reg_or_imm));

    // MUX for Reg2
    assign dealt_reg2 = (reg2_sel == 2'h0) ? result_MEM :
                                            ((reg2_sel == 2'h1) ? data_WB : reg2_EX);


    // // MUX for result (ALU or PC_EX)
    // assign result = load_npc_EX ? PC_EX : ALU_out;
    // MUX for result (ALU or PC_EX)  
    //TODO: CSR debug
    assign result = load_npc_EX ? PC_EX : (is_csr_out ? csr_read_data : ALU_out);


    //Module connections
    // ---------------------------------------------
    // PC-Generator
    // ---------------------------------------------


    NPC_Generator NPC_Generator1(
        .PC(PC_4),
        .jal_target(jal_target),
        .jalr_target(ALU_out),
        .br_target(br_target),
        .jal(jal),
        .jalr(jalr_EX),
        .br(br),
        .NPC(NPC),
        //Lab4
        .btb_if(btb_if),
        .btb_ex(btb_ex),
        .if_prediction_true(if_prediction_true),
        .prediction_if(prediction_if),
        .PC_EX(PC_EX),
        //Lab4 phase 2
        .bht_if(bht_if),
        .bht_ex(bht_ex)
    );


    PC_IF PC_IF1(
        .clk(CPU_CLK),
        .bubbleF(bubbleF),
        .flushF(flushF),
        .NPC(NPC),
        .PC(PC_IF)
    );



    // ---------------------------------------------
    // IF stage
    // ---------------------------------------------

    PC_ID PC_ID1(
        .clk(CPU_CLK),
        .bubbleD(bubbleD),
        .flushD(flushD),
        .PC_IF(PC_4),
        .PC_ID(PC_ID)
    );


    IR_ID IR_ID1(
        .clk(CPU_CLK),
        .bubbleD(bubbleD),
        .flushD(flushD),
        .write_en(|CPU_Debug_InstCache_WE2),
        .addr(PC_IF[31:2]),
        .debug_addr(CPU_Debug_InstCache_A2[31:2]),
        .debug_input(CPU_Debug_InstCache_WD2),
        .inst_ID(inst_ID),
        .debug_data(CPU_Debug_InstCache_RD2)
    );



    // ---------------------------------------------
    // ID stage
    // ---------------------------------------------


    RegisterFile RegisterFile1(
        .clk(CPU_CLK),
        .rst(CPU_RST),
        .write_en(reg_write_en_WB),
        .addr1(inst_ID[19:15]),
        .addr2(inst_ID[24:20]),
        .wb_addr(reg_dest_WB),
        .wb_data(data_WB),
        .reg1(reg1),
        .reg2(reg2)
    );

    ControllerDecoder ControllerDecoder1(
        .inst(inst_ID),
        .jal(jal),
        .jalr(jalr_ID),
        .op2_src(op2_src),
        .ALU_func(ALU_func_ID),
        .br_type(br_type_ID),
        .load_npc(load_npc_ID),
        .wb_select(wb_select_ID),
        .load_type(load_type_ID),
        .src_reg_en(src_reg_en_ID),
        .reg_write_en(reg_write_en_ID),
        .cache_write_en(cache_write_en_ID),
        .alu_src1(alu_src1_ID),
        .alu_src2(alu_src2_ID),
        .imm_type(imm_type),
    );

    ImmExtend ImmExtend1(
        .inst(inst_ID[31:7]),
        .imm_type(imm_type),
        .imm(imm)
    );


    PC_EX PC_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .PC_ID(PC_ID),
        .PC_EX(PC_EX)
    );

    BR_Target_EX BR_Target_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .address(jal_target),
        .address_EX(br_target)
    );

    Op1_EX Op1_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .reg1(reg1),
        .reg1_EX(reg1_EX)
    );

    Op2_EX Op2_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .op2(op2),
        .reg_or_imm(reg_or_imm)
    );

    Reg2_EX Reg2_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .reg2(reg2),
        .reg2_EX(reg2_EX)
    );

    Addr_EX Addr_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .reg1_src_ID(inst_ID[19:15]),
        .reg2_src_ID(inst_ID[24:20]),
        .reg_dest_ID(inst_ID[11:7]),
        .reg1_src_EX(reg1_src_EX),
        .reg2_src_EX(reg2_src_EX),
        .reg_dest_EX(reg_dest_EX)
    );


    wire [6:0] opcode_EX;
    Ctrl_EX Ctrl_EX1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .jalr_ID(jalr_ID),
        .ALU_func_ID(ALU_func_ID),
        .br_type_ID(br_type_ID),
        .load_npc_ID(load_npc_ID),
        .wb_select_ID(wb_select_ID),
        .load_type_ID(load_type_ID),
        .src_reg_en_ID(src_reg_en_ID),
        .reg_write_en_ID(reg_write_en_ID),
        .cache_write_en_ID(cache_write_en_ID),
        .alu_src1_ID(alu_src1_ID),
        .alu_src2_ID(alu_src2_ID),
        .jalr_EX(jalr_EX),
        .ALU_func_EX(ALU_func_EX),
        .br_type_EX(br_type_EX),
        .load_npc_EX(load_npc_EX),
        .wb_select_EX(wb_select_EX),
        .load_type_EX(load_type_EX),
        .src_reg_en_EX(src_reg_en_EX),
        .reg_write_en_EX(reg_write_en_EX),
        .cache_write_en_EX(cache_write_en_EX),
        .alu_src1_EX(alu_src1_EX),
        .alu_src2_EX(alu_src2_EX)
    );

    //TODO: CSR debug
    CSRAddrEx CsrAddrEx1(
        .clk(CPU_CLK),
        .bubbleE(bubbleE),
        .flushE(flushE),
        .csr_addr_in(inst_ID[31:20]),
        .csr_addr_out(csr_addr_EX),
        .func3_in(inst_ID[14:12]),
        .func3_out(csr_funct3_out),
        .zimm_in(inst_ID[19:15]),
        .zimm_out(csr_zimm_out),
        .csr_write_en_in(csr_write_en_in),
        .csr_write_en_out(csr_write_en_out),
        .is_csr_in(is_csr_in),
        .is_csr_out(is_csr_out)
    );

    // ---------------------------------------------
    // EX stage
    // ---------------------------------------------

    //TODO: CSR debug
    ControlAndStatusRegister csr(
        .clk(CPU_CLK),
        .rst(CPU_RST),
        .reg1(reg1_EX),
        .zimm(csr_zimm_out),
        .func3(csr_funct3_out),
        .read_reg_addr(csr_addr_EX),
        .csr_write_en(csr_write_en_out),
        .read_reg_data(csr_read_data),
        .is_csr(is_csr_out)
    );

    ALU ALU1(
        .op1(ALU_op1),
        .op2(ALU_op2),
        .ALU_func(ALU_func_EX),
        .ALU_out(ALU_out)
    );

    BranchDecision BranchDecision1(
        .reg1(ALU_op1),
        .reg2(dealt_reg2),
        .br_type(br_type_EX),
        .br(br)
    );


    Result_MEM Result_MEM1(
        .clk(CPU_CLK),
        .bubbleM(bubbleM),
        .flushM(flushM),
        .result(result),
        .result_MEM(result_MEM)
    );

    Reg2_MEM Reg2_MEM1(
        .clk(CPU_CLK),
        .bubbleM(bubbleM),
        .flushM(flushM),
        .reg2_EX(dealt_reg2),
        .reg2_MEM(reg2_MEM)
    );

    Addr_MEM Addr_MEM1(
        .clk(CPU_CLK),
        .bubbleM(bubbleM),
        .flushM(flushM),
        .reg_dest_EX(reg_dest_EX),
        .reg_dest_MEM(reg_dest_MEM)
    );



    Ctrl_MEM Ctrl_MEM1(
        .clk(CPU_CLK),
        .bubbleM(bubbleM),
        .flushM(flushM),
        .wb_select_EX(wb_select_EX),
        .load_type_EX(load_type_EX),
        .reg_write_en_EX(reg_write_en_EX),
        .cache_write_en_EX(cache_write_en_EX),
        .wb_select_MEM(wb_select_MEM),
        .load_type_MEM(load_type_MEM),
        .reg_write_en_MEM(reg_write_en_MEM),
        .cache_write_en_MEM(cache_write_en_MEM)
    );



    // ---------------------------------------------
    // MEM stage
    // ---------------------------------------------
    wire miss;
    assign debug_miss = miss;
    WB_Data_WB WB_Data_WB1(
        .clk(CPU_CLK),
        .bubbleW(bubbleW),
        .flushW(flushW),
        .wb_select(wb_select_MEM),
        .load_type(load_type_MEM),
        .write_en(cache_write_en_MEM),
        .debug_write_en(CPU_Debug_DataCache_WE2),
        .addr(result_MEM),
        .debug_addr(CPU_Debug_DataCache_A2),
        .in_data(reg2_MEM),
        .debug_in_data(CPU_Debug_DataCache_WD2),
        .debug_out_data(CPU_Debug_DataCache_RD2),
        .data_WB(data_WB),
        //Lab3
        .miss(miss),
        .rst(CPU_RST),
        .debug_cache_hit(debug_cache_hit),
        .total_count(total_count)
    );


    Addr_WB Addr_WB1(
        .clk(CPU_CLK),
        .bubbleW(bubbleW),
        .flushW(flushW),
        .reg_dest_MEM(reg_dest_MEM),
        .reg_dest_WB(reg_dest_WB)
    );

    Ctrl_WB Ctrl_WB1(
        .clk(CPU_CLK),
        .bubbleW(bubbleW),
        .flushW(flushW),
        .reg_write_en_MEM(reg_write_en_MEM),
        .reg_write_en_WB(reg_write_en_WB)
    );


    // ---------------------------------------------
    // WB stage
    // ---------------------------------------------



    // ---------------------------------------------
    // Harzard Unit
    // ---------------------------------------------
    HarzardUnit HarzardUnit1(
        .rst(CPU_RST),
        .reg1_srcD(inst_ID[19:15]),
        .reg2_srcD(inst_ID[24:20]),
        .reg1_srcE(reg1_src_EX),
        .reg2_srcE(reg2_src_EX),
        .reg_dstE(reg_dest_EX),
        .reg_dstM(reg_dest_MEM),
        .reg_dstW(reg_dest_WB),
        .br(br),
        .jalr(jalr_EX),
        .jal(jal),
        .src_reg_en(src_reg_en_EX),
        .wb_select(wb_select_EX),
        .reg_write_en_MEM(reg_write_en_MEM),
        .reg_write_en_WB(reg_write_en_WB),
        .alu_src1(alu_src1_EX),
        .alu_src2(alu_src2_EX),
        .flushF(flushF),
        .bubbleF(bubbleF),
        .flushD(flushD),
        .bubbleD(bubbleD),
        .flushE(flushE),
        .bubbleE(bubbleE),
        .flushM(flushM),
        .bubbleM(bubbleM),
        .flushW(flushW),
        .bubbleW(bubbleW),
        .op1_sel(op1_sel),
        .op2_sel(op2_sel),
        .reg2_sel(reg2_sel),
        //Lab3
        .miss(miss),
        //Lab4
        .btb_ex(btb_ex),
        .btb_operation(btb_operation),
        //Lab4
        .bht_ex(bht_ex),
        .if_prediction_true(if_prediction_true)
    );  
    	         
endmodule